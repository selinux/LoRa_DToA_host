seba@t440p.8504:1498739642